module IntructionFetch(output logic[31:0] encoded_value);

endmodule: InstructionFetch