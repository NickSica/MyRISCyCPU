// Code your testbench here
// or browse Examples
// https://github.com/RobertBaruch/lmarv/blob/master/lmarv-1/riscv-instructions-book/instr.pdf
// zipcpu.com/tutorial
// nandland.com