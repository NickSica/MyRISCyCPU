

module RAM
    (input logic clk,
    flags.src fsrc);
    

endmodule: RAM


