module Execute();

endmodule: Execute