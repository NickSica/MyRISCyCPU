

module ControlPath
    (input clk,
    flags.src fsrc);

    logic[4:0] prev_rd;
    
    

endmodule: ControlPath


