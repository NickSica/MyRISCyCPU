module Decode(input logic[31:0] encoded_value);

endmodule: Decode