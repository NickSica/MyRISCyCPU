module alu(input logic rd, input logic op1, input logic op2);
    
  
endmodule: alu